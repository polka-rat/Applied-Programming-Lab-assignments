.circuit
V1   1 GND  dc 2
R1   1   2     2
R2   2 GND     1
R3  2   1   2
.end
