.circuit
v1 1 GND dc 0
v2 GND 3 dc 15 
r1 1 2 10000 
r2 2 3 8100 
r3 2 GND 4700 
.end