Multiple dc sources 
.circuit
v1 1 GND dc 24
v2 3 GND dc 15
r1 1 2 10000
r2 2 3 8100
r3 2 GND 4700 
.end 